// chuanjun zhang
// 10111序列检测，要求非交叠检测（即对于101110111只检测到一次）；
// 使用三段式fsm实现；
// 寄存器输出且同步输出结果；
// 低电平复位；

// 总结：使用Moore状态机，状态数量 = 序列元素个数 + 1；
// 多的一个状态为idle mode（空闲模式：一种设备或系统在未执行任何任务时的状态，通常为了节省能源或等待新任务）；

module serial_10111_check(


);




module
